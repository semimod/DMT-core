HICUM2v2.40 Amplifier in Time Domain

vcc cc 0 1
vin b 0 ac 1 dc 0.94 sin 0.94 50m 700G
rl c cc 10
q1 c b 0 0 hicum_va

.temp 24
.control
option method=gear
set filetype=ascii
*set appendwrite
set wr_vecnames
set wr_singlescal
tran 0.001p 0.02n
wrdata output_tran all
.endc
.model hicum_va NPN level=8
*Transfer current
+ c10 = 9.074e-030
+ qp0 = 1.008e-013
+ ich = 0
+ hf0 = 40
+ hfe = 10.01
+ hfc = 20.04
+ hjei = 3.382
+ ahjei = 3
+ rhjei = 2
+ hjci = 0.2
*
*Base-Emitter diode currents
+ ibeis = 1.328e-019
+ mbei = 1.027
+ ireis = 1.5e-015
+ mrei = 2
+ ibeps = 1.26e-019
+ mbep = 1.042
+ ireps = 1.8e-015
+ mrep = 1.8
+ mcf = 1
*
*Transit time for excess recombination current at b-c barrier
+ tbhrec = 1e-010
*
*Base-Collector diode currents
+ ibcis = 4.603e-017
+ mbci = 1.15
+ ibcxs = 0
+ mbcx = 1
*
*Base-Emitter tunneling current
+ ibets = 0.02035
+ abet = 24
+ tunode = 1
*
*Base-Collector avalanche current
+ favl = 18.96
+ qavl = 5.092e-014
+ alfav = -0.0024
+ alqav = -0.0006284
+ kavl = 0.0
+ alkav = 0.0
*
*Series resistances
+ rbi0 = 4.444
+ rbx = 2.568
+ fgeo = 0.7409
+ fdqr0 = 0
+ fcrbi = 0
+ fqi = 1
+ re = 1.511
+ rcx = 2.483
*
*Substrate transistor
+ itss = 1.143e-017
+ msf = 1.056
+ iscs = 4.60106e-015
+ msc = 1.018
+ tsf = 0
*
*Intra-device substrate coupling
+ rsu = 500
+ csu = 6.4e-014
*
*Depletion Capacitances
+ cjei0 = 8.869e-015
+ vdei = 0.714
+ zei = 0.2489
+ ajei = 1.65
+ cjep0 = 2.178e-015
+ vdep = 0.8501
+ zep = 0.2632
+ ajep = 1.6
+ cjci0 = 3.58e-015
+ vdci = 0.8201
+ zci = 0.2857
+ vptci = 1.79
+ cjcx0 = 0
+ vdcx = 0.8201
+ zcx = 0.2863
+ vptcx = 1.977
+ fbcpar = 0.3
+ fbepar = 1
+ cjs0 = 2.6e-014
+ vds = 0.9997
+ zs = 0.4295
+ vpts = 100
+ cscp0 = 1.4e-014
+ vdsp = 0
+ zsp = 0.35
+ vptsp = 4
*
*Diffusion Capacitances
+ t0 = 2.089e-013
+ dt0h = 8e-014
+ tbvl = 8.25e-014
+ tef0 = 3.271e-013
+ gtfe = 3.548
+ thcs = 5.001e-012
+ ahc = 0.05
+ fthc = 0.7
+ rci0 = 9.523
+ vlim = 0.6999
+ vces = 0.01
+ vpt = 2
+ aick = 1e-3
+ delck = 2
+ tr = 0
+ vcbar = 0.04
+ icbar = 0.01
+ acbar = 1.5
*
*Isolation Capacitances
+ cbepar = 0
+ cbcpar = 0
*
*Non-quasi-static Effect
+ flnqs = 1
+ alqf = 1
+ alit = 1
*
*Noise
+ kf = .3e-16
+ af = .75
+ cfbe = -1
+ flcono = 0
+ kfre = 0.0
+ afre = 2.0
*
*Lateral Geometry Scaling (at high current densities)
+ latb = 0.0
+ latl = 0.0
*
*Temperature dependence
+ vgb = 0.91
+ alt0 = 0.004
+ kt0 = 6.588e-005
+ zetaci = 0.58
+ alvs = 0.001
+ alces = -0.2286
+ zetarbi = 0.3002
+ zetarbx = 0.06011
+ zetarcx = -0.02768
+ zetare = -0.9605
+ zetacx = 0
+ vge = 1.17
+ vgc = 1.17
+ vgs = 1.049
+ f1vg = -0.000102377
+ f2vg = 0.00043215
+ zetact = 5
+ zetabet = 4.892
+ alb = 0
+ dvgbe = 0
+ zetahjei = -0.5
+ zetavgbe = 0.7
*
*Self-Heating
+ flsh = 0
+ rth = 1113.4
+ cth = 6.841e-012
+ zetarth = 0
+ alrth = 0.002
*
*Compatibility with V2.1
+ flcomp = 2.3
*
*Circuit simulator specific parameters
+ tnom = 26.85
*+ dt = 0

.end
